package g_inverter_tb_parampkg;
  parameter Latency = 41;
  parameter Input_Width = 104;
  parameter Input_Ports = 250;
  parameter Enable_Port = 0;
  parameter Logical_Function = AND;
endpackage

package g_addshiftreg_tb_parampkg;
  parameter Latency = 56;
  parameter Width = 246;
  parameter Enable_Port = 1;
endpackage

package g_simpledpram_tb_parampkg;
  parameter RAM_WIDTH = 206;
  parameter RAM_DEPTH = 61264;
  parameter INIT_FILE = "All zeros";
  parameter Write_Mode = 0;
  parameter Enable_Port_A = 0;
  parameter Reset_Port_A = 0;
  parameter Enable_Port_B = 1;
  parameter Reset_Port_B = 1;
  parameter Two_CLK = 0;
  parameter Latency = 1;
endpackage

package g_cmultrom_tb_parampkg;
  parameter Latency = 154;
  parameter Width = 29;
  parameter Enable_Port = 1;
  parameter Signed_Unsigned = 0;
  parameter Constant_Value = 250;
  parameter DATA_FILE = "C:\\questasim64_10.4c\\examples\\cmultromtables\\g_cmultrom_data_250.txt";
endpackage

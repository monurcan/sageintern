package g_relational_tb_parampkg;
  parameter Latency = 187;
  parameter Input_Width = 68;
  parameter Signed_Unsigned = 0;
  parameter Enable_Port = 0;
  parameter Comparison = "A>=B";
endpackage

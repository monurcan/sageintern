package g_fifo_tb_parampkg;
  parameter FIFO_WIDTH = 77;
  parameter FIFO_DEPTH = 44994;
  parameter FWFT = 0;
  parameter Enable_Port = 0;
  parameter Reset_Port = 1;
  parameter Data_Count_Port = 1;
  parameter Almost_Empty_Port = 0;
  parameter Almost_Full_Port = 1;
  parameter Almost_Empty_Treshold = 20983;
  parameter Almost_Full_Treshold = 22866;
endpackage

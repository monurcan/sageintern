package g_accumulator_tb_parampkg;
  parameter Operation = 0;
  parameter Latency = 10;
  parameter Signed_Unsigned = 0;
  parameter Width = 4;
  parameter Reset_Port = 1;
  parameter Reset_Bypass = 0;
  parameter Enable_Port = 0;
endpackage

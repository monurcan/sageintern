package g_mux_tb_parampkg;
  parameter Latency = 98;
  parameter Input_Width = 192;
  parameter Input_Ports = 186;
  parameter Enable_Port = 1;
endpackage

package g_rom_tb_parampkg;
  parameter Latency = 239;
  parameter Width = 174;
  parameter Depth = 53656;
  parameter Enable_Port = 0;
  parameter DATA_FILE = "C:\\questasim64_10.4c\\examples\\g_rom_data.txt";
endpackage

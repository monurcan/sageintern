package g_addsub_tb_parampkg;
  parameter Operation = 2;
  parameter Latency = 44;
  parameter Signed_Unsigned = 1;
  parameter Width = 105;
  parameter Reset_Port = 0;
  parameter Carry_In_Port = 0;
  parameter Carry_Out_Port = 1;
  parameter Enable_Port = 0;
endpackage

package g_spram_tb_parampkg;
  parameter RAM_WIDTH = 64;
  parameter RAM_DEPTH = 5823;
  parameter INIT_FILE = "All zeros";
  parameter Memory_Type = 1;
  parameter Write_Mode = 0;
  parameter Enable_Port = 1;
  parameter Reset_Port = 1;
  parameter Latency = 132;
endpackage

package g_treshold_tb_parampkg;
  parameter Latency = 100;
  parameter Port_Width = 5;
  parameter Enable_Port = 1;
endpackage

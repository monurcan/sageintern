package g_register_tb_parampkg;
  parameter Initial_Value = 1579;
  parameter Width = 99;
  parameter Enable_Port = 0;
  parameter Reset_Port = 1;
endpackage

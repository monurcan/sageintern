package g_leadingdet_tb_parampkg;
  parameter A_Width = 215;
  parameter Latency = 47;
  parameter Detect_from = 1;
  parameter Detect_Value = 1;
  parameter Enable_Port = 0;
endpackage

package g_multiplierus_tb_parampkg;
  parameter A_Width = 79;
  parameter B_Width = 204;
  parameter Enable_Port = 0;
endpackage

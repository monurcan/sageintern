package g_constant_tb_parampkg;
  parameter Constant_Value = -1043810061;
  parameter Port_Width = 201;
endpackage

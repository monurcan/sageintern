package g_slice_tb_parampkg;
  parameter Input_Width = 172;
  parameter Slice_Width = 125;
  parameter Specify_range_as = 3;
  parameter High_Bit = 155;
  parameter Low_Bit = 31;
endpackage

package g_cmultlut_tb_parampkg;
  parameter Latency = 150;
  parameter Signed_Unsigned = 0;
  parameter A_Width = 65;
  parameter Constant_Value = 201;
  parameter Enable_Port = 0;
  parameter Reset_Port = 0;
endpackage

package g_multiplier_tb_parampkg;
  parameter Latency = 254;
  parameter Signed_Unsigned = 0;
  parameter A_Width = 19;
  parameter B_Width = 207;
  parameter Enable_Port = 0;
endpackage

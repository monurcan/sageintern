package g_counter_tb_parampkg;
  parameter Count_Limit = 252;
  parameter Width = 235;
  parameter Direction = 2;
  parameter G_Initial_Value = 246;
  parameter Step = 155;
  parameter Out_type = 1;
  parameter Reset_Port = 1;
  parameter Load_Port = 1;
  parameter Enable_Port = 1;
  parameter Free_or_Limited = 0;
endpackage

package g_delay_tb_parampkg;
  parameter Latency = 226;
  parameter Width = 72;
  parameter Reset_Port = 1;
  parameter Enable_Port = 1;
endpackage

package g_truedpram_tb_parampkg;
  parameter RAM_WIDTH = 169;
  parameter RAM_DEPTH = 18786;
  parameter INIT_FILE = "All zeros";
  parameter Write_Mode = 0;
  parameter Enable_Port_A = 0;
  parameter Reset_Port_A = 1;
  parameter Enable_Port_B = 0;
  parameter Reset_Port_B = 0;
  parameter Two_CLK = 1;
  parameter Latency_A = 13;
  parameter Latency_B = 1;
endpackage

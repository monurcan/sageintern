package g_logical_tb_parampkg0;
  parameter Latency = 60;
  parameter Input_Width = 75;
  parameter Input_Ports = 22;
  parameter Enable_Port = 1;
  parameter Logical_Function = "XOR";
endpackage
package g_logical_tb_parampkg1;
  parameter Latency = 76;
  parameter Input_Width = 30;
  parameter Input_Ports = 201;
  parameter Enable_Port = 0;
  parameter Logical_Function = "INVALID";
endpackage
package g_logical_tb_parampkg2;
  parameter Latency = 181;
  parameter Input_Width = 103;
  parameter Input_Ports = 409;
  parameter Enable_Port = 1;
  parameter Logical_Function = "XNOR";
endpackage
package g_logical_tb_parampkg3;
  parameter Latency = 129;
  parameter Input_Width = 18;
  parameter Input_Ports = 163;
  parameter Enable_Port = 1;
  parameter Logical_Function = "NAND";
endpackage
package g_logical_tb_parampkg4;
  parameter Latency = 243;
  parameter Input_Width = 62;
  parameter Input_Ports = 173;
  parameter Enable_Port = 0;
  parameter Logical_Function = "INVALID";
endpackage

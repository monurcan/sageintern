package g_barrelshift_tb_parampkg;
  parameter Latency = 165;
  parameter A_Width = 85;
  parameter Direction = 5;
  parameter Enable_Port = 1;
endpackage
